class uvm_template_env extends uvm_env;


endclass : uvm_template_env