package uvm_template_env_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import uvm_template_seq_pkg::*;
  import uvm_template_agent_pkg::*;
  `include "uvm_template_sb.sv"
  `include "uvm_template_env.sv"

endpackage : uvm_template_env_pkg
