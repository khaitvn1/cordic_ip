package uvm_template_test_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import uvm_template_env_pkg::*;
  import uvm_template_seq_pkg::*;
  `include "uvm_template_base_test.svh"
  `include "uvm_template_test_lib.sv"
  
endpackage : uvm_template_test_pkg
