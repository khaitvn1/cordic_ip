class base_cordic_seq extends uvm_sequence #(cordic_seq_item);

endclass : base_cordic_seq