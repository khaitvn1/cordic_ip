class simple_cordic_test extends base_cordic_test;

endclass : simple_cordic_test
