class base_uvm_template_seq extends uvm_sequence #(uvm_template_seq_item);

endclass : base_uvm_template_seq