class cordic_agent extends uvm_agent;

endclass : cordic_agent