class uvm_template_seq_item extends uvm_sequence_item;


endclass : uvm_template_seq_item