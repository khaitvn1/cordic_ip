package uvm_template_agent_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import uvm_template_seq_pkg::*;
    `include "uvm_template_monitor.sv"
    `include "uvm_template_driver.sv"
    `include "uvm_template_sequencer.sv"
    `include "uvm_template_agent.sv"
endpackage : uvm_template_agent_pkg