class cordic_sb extends uvm_scoreboard;

endclass : cordic_sb
