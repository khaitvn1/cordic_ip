class uvm_template_monitor extends uvm_monitor;


endclass : uvm_template_monitor