class cordic_seq_item extends uvm_sequence_item;


endclass : cordic_seq_item