class uvm_template_agent extends uvm_agent;

endclass : uvm_template_agent