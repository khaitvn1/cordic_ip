class simple_cordic_seq extends base_cordic_seq;

endclass : simple_cordic_seq