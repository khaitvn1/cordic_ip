class cordic_env extends uvm_env;


endclass : cordic_env