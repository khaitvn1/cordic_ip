class cordic_monitor extends uvm_monitor;


endclass : cordic_monitor