package cordic_seq_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import cordic_tb_pkg::*;
    import cordic_pkg::*;
    `include "cordic_seq_item.sv"
    `include "cordic_sequence.svh"
    `include "cordic_seq_lib.sv"
endpackage : cordic_seq_pkg
