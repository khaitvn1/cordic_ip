class cordic_driver extends uvm_driver #(cordic_seq_item);

endclass : cordic_driver