class uvm_template_sequencer extends uvm_sequencer #(uvm_template_seq_item);


endclass : uvm_template_sequencer