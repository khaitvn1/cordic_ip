class base_cordic_test extends uvm_test;

endclass : base_cordic_test