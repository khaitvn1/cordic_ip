package uvm_template_seq_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "uvm_template_seq_item.sv"
  `include "uvm_template_sequence.svh"
  `include "uvm_template_seq_lib.sv"
  
endpackage : uvm_template_seq_pkg
