package cordic_test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    import cordic_tb_pkg::*;
    import cordic_pkg::*;
    import cordic_env_pkg::*;
    import cordic_seq_pkg::*;
    `include "cordic_base_test.svh"
    `include "cordic_test_lib.sv"
endpackage : cordic_test_pkg
