class base_uvm_template_test extends uvm_test;

endclass : base_uvm_template_test