class uvm_template_sb extends uvm_scoreboard;

endclass : uvm_template_sb
