class cordic_sequencer extends uvm_sequencer #(cordic_seq_item);


endclass : cordic_sequencer