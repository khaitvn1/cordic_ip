class uvm_template_driver extends uvm_driver #(uvm_template_seq_item);

endclass : uvm_template_driver